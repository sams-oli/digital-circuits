`ifndef ALUOP
`define ALUOP

`define ALU_ADDU 4'd0
`define ALU_SUBU 4'd1
`define ALU_SLT  4'd2
`define ALU_SLTU 4'd3
`define ALU_AND  4'd4
`define ALU_OR   4'd5
`define ALU_XOR  4'd6
`define ALU_LUI  4'd7
`define ALU_SLL  4'd8
`define ALU_SRL  4'd9
`define ALU_SRA  4'd10
`define ALU_NOR  4'd11
`define ALU_XXX  4'd15

`endif // ALUOP
