// Module Purpose:
//		Este módulo provê uma saída de único ciclo, baseada em um push button
// -----------------------------------------------------------------------------
//	Params:		Este módulo não é parametrizado.
//	Inputs:		Ver documento do laboratório.
//	Outputs:		Ver documento do laboratório.
// -----------------------------------------------------------------------------
module level2pulse (
	//------------------------------------------------------------------
	//	Entradas Clock & Reset
	//------------------------------------------------------------------
	input wire clock,
	input wire reset,
	//------------------------------------------------------------------
	
	//------------------------------------------------------------------
	//	Entradas
	//------------------------------------------------------------------
	input wire level,
	//------------------------------------------------------------------
	
	//------------------------------------------------------------------
	//	Saídas
	//------------------------------------------------------------------
	output logic pulse
	//------------------------------------------------------------------
);

	//--------------------------------------------------------------------------
	//	Codificação dos estados
	//--------------------------------------------------------------------------
	
	parameter [3:0] E0  = 4'b0000,
                  	E1 = 4'b0001,
                  	E2 = 4'b0010;
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Declaração dos wires
	//--------------------------------------------------------------------------
	
	reg [3:0] state, prox;
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Lógica
	//--------------------------------------------------------------------------
	
	always @(posedge clock or negedge reset)
    	if (!reset) state <= E0;
    	else        state <= prox;

	always @(state or level) begin
   		prox = 4'bx;
    	pulse = 1'b0;

    case (state)
      E0 :   if (!level)       	prox = E1;
             else           	prox = E0;

      E1: begin
               	pulse = 1'b1;
				prox = E2;
	end

      E2:   if (!level)      prox = E2;
            else           prox = E0;

    endcase
end

	//--------------------------------------------------------------------------
endmodule // level2pulse
